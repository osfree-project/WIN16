# Translation by Martin Str�mberg <ams@ludd.luth.se>.
0.0:Visa inneh�llet i en textfil en sk�rm i taget
0.1:Anv�ndning
0.2:kommando
0.3:fil
0.4:Tillg�ngliga tangenter
0.5:Nn
0.6:N�sta fil
0.7:Qq
0.8:Avsluta program
0.9:Mellanslag
0.10:N�sta sida
1.0:Ok�nd option
1.1:Ingen s�dan fil
1.2:Kan inte �ppna filen
2.0:Mera
2.1:<STDIN>
